
module top_level(
    input clk,
    input clk_en,
    input sync_rst
);



endmodule
